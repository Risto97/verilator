module t(
);
    if(1) begin : block1 
        assign wire_l1 = wire_l0;
        wire wire_l1;
    end

    wire wire_l0;
endmodule

